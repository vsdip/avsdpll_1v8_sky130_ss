* SPICE3 file created from CP.ext - technology: sky130A
.include ~/Characterization-TCL-flow-for-8x-PLL-Clock-Multiplier-for-sky130-Process-Corners/sky130nm.lib
.option scale=0.01u

*.subckt CP VDD GND Up Down Out ENb
XM1000 a_86_73# a_125_486# a_248_475# VDD sky130_fd_pr__pfet_01v8 w=1800 l=15
+  ad=68834 pd=4394 as=62586 ps=3832
XM1001 GND a_340_202# a_462_191# GND sky130_fd_pr__nfet_01v8 w=480 l=15
+  ad=20982 pd=1602 as=23046 ps=1312
XM1002 a_86_73# a_125_486# a_125_486# VDD sky130_fd_pr__pfet_01v8 w=44 l=15
+  ad=0 pd=0 as=1452 ps=154
XM1003 a_248_475# a_134_73# Out VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=0 pd=0 as=1386 ps=150
XM1004 a_134_73# Down GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1188 pd=138 as=0 ps=0
XM1005 a_248_475# Down a_248_427# VDD sky130_fd_pr__pfet_01v8 w=540 l=15
+  ad=0 pd=0 as=17820 ps=1146
XM1006 a_258_74# Up GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1188 pd=138 as=0 ps=0
XM1007 GND a_340_202# a_340_202# GND sky130_fd_pr__nfet_01v8 w=44 l=15
+  ad=0 pd=0 as=1452 ps=154
XM1008 a_462_143# a_462_143# a_86_73# VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1386 pd=150 as=0 ps=0
XM1009 Out Up a_462_191# GND sky130_fd_pr__nfet_01v8 w=42 l=15
+  ad=1386 pd=150 as=0 ps=0
XM1010 a_248_427# a_248_427# GND GND sky130_fd_pr__nfet_01v8 w=42 l=15
+  ad=1386 pd=150 as=0 ps=0
XM1011 VDD ENb a_86_73# VDD sky130_fd_pr__pfet_01v8 w=1800 l=15
+  ad=50400 pd=3656 as=0 ps=0
XM1012 a_462_191# a_258_74# a_462_143# GND sky130_fd_pr__nfet_01v8 w=540 l=15
+  ad=0 pd=0 as=17820 ps=1146
XM1013 a_258_74# Up a_86_73# VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=2376 pd=210 as=0 ps=0
XM1014 a_134_73# Down a_86_73# VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=2376 pd=210 as=0 ps=0
C0 a_258_74# VDD 0.08fF
C1 VDD a_248_475# 1.36fF
C2 a_125_486# VDD 0.05fF
C3 Up a_462_143# 0.08fF
C4 a_134_73# a_86_73# 0.21fF
C5 Out a_248_475# 0.40fF
C6 a_86_73# a_462_191# 0.01fF
C7 VDD a_86_73# 5.67fF
C8 VDD a_134_73# 0.04fF
C9 a_248_427# Down 0.00fF
C10 Up a_340_202# 0.02fF
C11 VDD a_462_191# 0.13fF
C12 a_258_74# a_462_143# 0.02fF
C13 Out a_86_73# 0.33fF
C14 a_258_74# a_248_427# 0.00fF
C15 a_248_427# a_248_475# 0.58fF
C16 Out a_134_73# 0.05fF
C17 Out a_462_191# 0.04fF
C18 Out VDD 1.46fF
C19 Up Down 0.14fF
C20 a_462_143# a_86_73# 0.16fF
C21 a_258_74# a_340_202# 0.13fF
C22 a_248_427# a_86_73# 0.25fF
C23 a_248_427# a_134_73# 0.09fF
C24 Up a_258_74# 0.08fF
C25 a_462_143# a_462_191# 0.72fF
C26 VDD a_462_143# 0.20fF
C27 a_248_427# a_462_191# 0.02fF
C28 VDD a_248_427# 0.17fF
C29 ENb Down 0.01fF
C30 a_134_73# a_340_202# 0.00fF
C31 a_258_74# Down 0.00fF
C32 Out a_462_143# 0.02fF
C33 Up a_86_73# 1.58fF
C34 a_125_486# Down 0.02fF
C35 Up a_134_73# 0.41fF
C36 a_340_202# a_462_191# 0.01fF
C37 ENb a_248_475# 0.00fF
C38 Out a_248_427# 0.00fF
C39 VDD a_340_202# 0.02fF
C40 a_125_486# ENb 0.10fF
C41 Up a_462_191# 0.09fF
C42 a_125_486# a_248_475# 0.02fF
C43 Up VDD 0.08fF
C44 a_86_73# Down 0.06fF
C45 a_134_73# Down 0.12fF
C46 a_248_427# a_462_143# 0.01fF
C47 a_258_74# a_86_73# 0.15fF
C48 a_248_475# a_86_73# 2.08fF
C49 VDD Down 0.03fF
C50 Out Up 0.03fF
C51 a_258_74# a_134_73# 0.05fF
C52 a_248_475# a_134_73# 0.02fF
C53 a_125_486# a_86_73# 0.06fF
C54 VDD ENb 0.16fF
C55 a_258_74# a_462_191# 0.00fF
C56 Up 0 0.07fF
C57 Out 0 2.98fF
C58 VDD 0 0.32fF
C59 a_462_143# 0 0.55fF
C60 a_462_191# 0 0.58fF
C61 a_340_202# 0 0.31fF
C62 a_258_74# 0 0.51fF
C63 a_134_73# 0 2.42fF
C64 a_248_427# 0 0.69fF
C65 a_248_475# 0 0.49fF
C66 a_125_486# 0 0.24fF
C67 a_86_73# 0 1.79fF


c90 Out GND 6fF
v1 VDD GND 1.8
*Up signal
v2 Up GND PULSE 0 1.8 4ns 6p 6p 100n 200n
v3 Down GND 0 
v4 ENb GND 0

.ic v(Out) = 0
.control
tran 1n 5u
plot v(Up) v(Down) v(Out)+2
.endc
