VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO FD
  CLASS CORE ;
  FOREIGN FD ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.350 BY 3.200 ;
  SITE unithddb1 ;
  PIN Clk_Out
    ANTENNADIFFAREA 0.318700 ;
    PORT
      LAYER li1 ;
        RECT 8.910 2.550 9.090 2.590 ;
        RECT 8.910 1.810 9.200 2.550 ;
        RECT 8.950 1.640 9.200 1.810 ;
        RECT 9.030 0.980 9.200 1.640 ;
        RECT 8.900 0.620 9.200 0.980 ;
    END
  END Clk_Out
  PIN GND
    ANTENNADIFFAREA 1.261200 ;
    PORT
      LAYER li1 ;
        RECT 0.410 0.320 0.580 1.110 ;
        RECT 1.520 0.320 1.690 1.110 ;
        RECT 4.250 0.320 4.420 1.100 ;
        RECT 6.910 0.320 7.080 1.110 ;
        RECT 8.420 0.320 8.640 0.910 ;
        RECT 0.000 0.150 9.350 0.320 ;
      LAYER mcon ;
        RECT 0.160 0.150 0.330 0.320 ;
        RECT 1.000 0.150 1.170 0.320 ;
        RECT 1.800 0.150 1.970 0.320 ;
        RECT 3.150 0.150 3.320 0.320 ;
        RECT 4.070 0.150 4.240 0.320 ;
        RECT 5.130 0.150 5.300 0.320 ;
        RECT 5.970 0.150 6.140 0.320 ;
        RECT 7.150 0.150 7.320 0.320 ;
        RECT 7.990 0.150 8.160 0.320 ;
        RECT 8.830 0.150 9.000 0.320 ;
      LAYER met1 ;
        RECT 0.000 0.000 9.350 0.480 ;
    END
  END GND
  PIN Clk_In
    ANTENNAGATEAREA 0.351000 ;
    PORT
      LAYER li1 ;
        RECT 6.490 2.160 6.660 2.500 ;
        RECT 0.000 1.310 0.660 1.480 ;
        RECT 2.370 0.740 2.700 0.920 ;
      LAYER mcon ;
        RECT 6.490 2.240 6.660 2.410 ;
        RECT 0.410 1.310 0.580 1.480 ;
        RECT 2.450 0.750 2.620 0.920 ;
      LAYER met1 ;
        RECT 0.350 2.180 1.570 2.500 ;
        RECT 6.440 2.490 6.720 2.500 ;
        RECT 0.350 1.270 0.640 2.180 ;
        RECT 1.320 2.070 1.570 2.180 ;
        RECT 6.430 2.070 6.720 2.490 ;
        RECT 1.320 1.820 6.720 2.070 ;
        RECT 0.360 0.980 0.640 1.270 ;
        RECT 0.360 0.690 2.710 0.980 ;
    END
  END Clk_In
  PIN VDD
    ANTENNADIFFAREA 1.829700 ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.830 9.320 3.020 ;
        RECT 0.410 1.730 0.580 2.830 ;
        RECT 1.520 1.730 1.690 2.830 ;
        RECT 4.250 1.720 4.420 2.830 ;
        RECT 6.910 1.730 7.080 2.830 ;
        RECT 8.410 2.220 8.640 2.830 ;
      LAYER mcon ;
        RECT 0.550 2.830 0.740 3.020 ;
        RECT 1.370 2.830 1.560 3.020 ;
        RECT 2.820 2.830 3.010 3.020 ;
        RECT 3.600 2.830 3.790 3.020 ;
        RECT 4.540 2.830 4.730 3.020 ;
        RECT 5.620 2.830 5.810 3.020 ;
        RECT 6.820 2.830 7.010 3.020 ;
        RECT 7.680 2.830 7.870 3.020 ;
        RECT 8.540 2.830 8.730 3.020 ;
      LAYER met1 ;
        RECT 0.000 2.720 9.320 3.200 ;
    END
  END VDD
  OBS
      LAYER li1 ;
        RECT 0.850 1.560 1.020 2.450 ;
        RECT 1.960 1.570 2.130 2.450 ;
        RECT 2.440 2.220 2.610 2.550 ;
        RECT 2.940 1.930 3.110 2.460 ;
        RECT 2.390 1.630 3.110 1.930 ;
        RECT 2.390 1.570 2.640 1.630 ;
        RECT 0.850 1.260 1.150 1.560 ;
        RECT 1.430 1.310 1.770 1.480 ;
        RECT 1.960 1.270 2.640 1.570 ;
        RECT 0.850 0.750 1.020 1.260 ;
        RECT 1.960 0.750 2.130 1.270 ;
        RECT 2.940 0.830 3.110 1.630 ;
        RECT 3.380 1.900 3.550 2.460 ;
        RECT 3.380 1.630 4.080 1.900 ;
        RECT 3.380 0.830 3.550 1.630 ;
        RECT 3.910 1.540 4.080 1.630 ;
        RECT 4.690 1.560 4.860 2.440 ;
        RECT 5.590 1.910 5.760 2.450 ;
        RECT 5.090 1.620 5.760 1.910 ;
        RECT 5.090 1.560 5.370 1.620 ;
        RECT 3.910 1.520 4.120 1.540 ;
        RECT 3.910 1.470 4.460 1.520 ;
        RECT 3.910 1.300 4.500 1.470 ;
        RECT 3.910 1.270 4.460 1.300 ;
        RECT 4.690 1.270 5.370 1.560 ;
        RECT 4.690 0.740 4.860 1.270 ;
        RECT 5.090 0.710 5.420 0.880 ;
        RECT 5.590 0.820 5.760 1.620 ;
        RECT 6.030 1.880 6.200 2.450 ;
        RECT 6.030 1.630 6.570 1.880 ;
        RECT 6.030 0.820 6.200 1.630 ;
        RECT 6.380 1.520 6.570 1.630 ;
        RECT 7.350 1.560 7.520 2.450 ;
        RECT 7.900 2.010 8.120 2.590 ;
        RECT 7.900 1.840 8.740 2.010 ;
        RECT 8.550 1.640 8.740 1.840 ;
        RECT 6.790 1.520 7.120 1.530 ;
        RECT 6.380 1.480 7.120 1.520 ;
        RECT 6.380 1.310 7.160 1.480 ;
        RECT 6.380 1.280 7.120 1.310 ;
        RECT 6.380 1.010 6.570 1.280 ;
        RECT 7.350 1.260 7.690 1.560 ;
        RECT 8.010 1.420 8.350 1.590 ;
        RECT 8.550 1.350 8.770 1.640 ;
        RECT 8.540 1.300 8.770 1.350 ;
        RECT 6.380 0.700 6.660 1.010 ;
        RECT 7.350 0.750 7.520 1.260 ;
        RECT 8.540 1.250 8.720 1.300 ;
        RECT 7.890 1.080 8.720 1.250 ;
        RECT 7.890 0.620 8.110 1.080 ;
      LAYER mcon ;
        RECT 2.440 2.290 2.610 2.470 ;
        RECT 0.910 1.320 1.080 1.490 ;
        RECT 1.520 1.310 1.690 1.480 ;
        RECT 5.170 0.710 5.340 0.880 ;
        RECT 7.440 1.320 7.610 1.490 ;
        RECT 8.100 1.420 8.270 1.590 ;
        RECT 6.460 0.770 6.630 0.940 ;
      LAYER met1 ;
        RECT 2.370 2.220 2.690 2.540 ;
        RECT 0.830 1.240 1.180 1.590 ;
        RECT 1.460 1.260 7.690 1.540 ;
        RECT 8.040 1.370 8.350 1.650 ;
        RECT 8.070 1.000 8.340 1.370 ;
        RECT 5.080 0.630 5.410 0.960 ;
        RECT 6.400 0.730 8.340 1.000 ;
        RECT 6.400 0.710 6.720 0.730 ;
        RECT 6.410 0.700 6.720 0.710 ;
      LAYER via ;
        RECT 2.400 2.250 2.660 2.510 ;
        RECT 0.880 1.290 1.140 1.550 ;
        RECT 5.110 0.660 5.380 0.930 ;
      LAYER met2 ;
        RECT 0.850 1.590 1.180 1.660 ;
        RECT 0.830 1.570 1.180 1.590 ;
        RECT 2.370 1.570 2.690 2.510 ;
        RECT 0.830 1.280 5.400 1.570 ;
        RECT 0.830 1.240 1.180 1.280 ;
        RECT 5.070 0.930 5.400 1.280 ;
        RECT 5.070 0.870 5.410 0.930 ;
        RECT 5.080 0.630 5.410 0.870 ;
  END
END FD
END LIBRARY

